module not_gate(input a, output b);
  assign b = ~a;
endmodule
